module build3;
endmodule
