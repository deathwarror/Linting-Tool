module forLoop(
  input wire in,
  output reg out);
  reg i[5];
  
  for( ;;)begin
    
  end
  
endmodule
