library verilog;
use verilog.vl_types.all;
entity Vending_Machine_TB is
end Vending_Machine_TB;
