library verilog;
use verilog.vl_types.all;
entity FlipFlops_TB is
end FlipFlops_TB;
