module assng(
  input wire bob,
  input wire boob,
  output reg tom
  );
  wire toon;
  assign toon = bob;
  assign toon=boob ;
  
  
endmodule
