module LineNum(
  input wire bob,
  output reg tom
  );
  
  parameter param = 1;
  
  wire one;
  reg two;
  
  always@(bob 
  or one)begin
    tom = bob;
  end
  
  assign one = two;
  
endmodule
