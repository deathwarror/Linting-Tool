module submod(
  input wire in,
  output reg out
  );
  radix rad_man(.in(in), . out ( out ) );
  
  
endmodule
