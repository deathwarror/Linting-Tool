library verilog;
use verilog.vl_types.all;
entity Sequence_Analyzer_TB is
end Sequence_Analyzer_TB;
