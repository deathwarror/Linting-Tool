library verilog;
use verilog.vl_types.all;
entity shell is
    port(
        bob             : in     vl_logic;
        bobby           : out    vl_logic
    );
end shell;
