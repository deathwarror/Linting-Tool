library verilog;
use verilog.vl_types.all;
entity Double_Sensitive_Clock_TB is
end Double_Sensitive_Clock_TB;
