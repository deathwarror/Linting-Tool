module Single_Assigned_Output(input wire a,b,c, output wire out);
  assign out = a+b+c;
endmodule
