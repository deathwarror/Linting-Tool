//this is a comment
module 
shell
(
input
 bob
 , 
 output
  bobby
  )
  ;
  // bob bbop
  /* oh no
  bob
  charsl*/
  reg tom;
//  input wire tommy;
endmodule
