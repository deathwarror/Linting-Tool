module build2 (a,b,c,d);
  input a, b, c;
  output wire d;
  wire e;
endmodule
