module param(
  input wire one,
  output reg two
  );
  
  parameter three = 5;
  localparam four = 6;

  parameter bob = three-1;
  parameter sue = bob-1;
  
endmodule
