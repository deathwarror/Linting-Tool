`default_nettype none
module build (
input wire f, g, a, b,c, 
input dd, input reg e,
output wire ch,
 wire bob);
//  assign ch = a+f;
  output bob;

  reg carla;
  reg bobby, bomber;
endmodule
